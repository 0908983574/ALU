module ALU   ( //Change what do you do verilog file ok i choose incomming change
    out, in
);
    input in;
    output out;

    assign out = in;
    assign out = in;
    
endmodule
