module ALU   ( //Change I don no verilog file
    out, in
);
    input in;
    output out;

    assign out = in;
    assign out = in;
    
endmodule
