module ALU   ( //Change verilog file
    out, in
);
    input in;
    output out;

    assign out = in;
    assign out = in;
    
endmodule
